module datapath (
    part,
    clock,
    value,
    positive,
    reset,
    counter,
    result
);

    input part;
    input clock;
    input [15:0] value;
    input positive;
    input reset;
    output [15:0] counter;
    output [15:0] result;

    /* signal declarations */
    wire [15:0] _65 = 16'b0000000000000000;
    wire [15:0] _64 = 16'b0000000000000000;
    wire _102;
    wire _100;
    wire _101;
    wire _103;
    wire [15:0] _104;
    wire _96;
    wire _92;
    wire _93;
    wire _90;
    wire _91;
    wire _94;
    wire _95;
    wire _97;
    wire [15:0] _98;
    wire _86;
    wire _84;
    wire _81;
    wire _82;
    wire _79;
    wire _80;
    wire _83;
    wire _85;
    wire _87;
    wire [15:0] _88;
    wire [41:0] _73 = 42'b000000000000000000000010100011110101110001;
    wire [25:0] _71 = 26'b00000000000000000000000000;
    wire [41:0] _72;
    wire [83:0] _74;
    wire [57:0] _75;
    wire [25:0] _70 = 26'b00000000000000000000000000;
    wire [83:0] _76;
    wire [15:0] _77;
    wire [15:0] _78;
    wire [15:0] _89;
    wire [15:0] _99;
    wire [15:0] _105;
    wire [15:0] _67 = 16'b0000000000000001;
    wire [15:0] _68;
    wire [15:0] _62 = 16'b0000000000000000;
    wire [15:0] _58 = 16'b0000000001100100;
    wire [41:0] _53 = 42'b000000000000000000000010100011110101110001;
    wire [25:0] _51 = 26'b00000000000000000000000000;
    wire [41:0] _52;
    wire [83:0] _54;
    wire [57:0] _55;
    wire [25:0] _50 = 26'b00000000000000000000000000;
    wire [83:0] _56;
    wire [15:0] _57;
    wire [31:0] _59;
    wire [15:0] _60;
    wire [15:0] _48 = 16'b0000000000110010;
    wire [15:0] _44 = 16'b0000000001100100;
    wire [41:0] _39 = 42'b000000000000000000000010100011110101110001;
    wire [25:0] _37 = 26'b00000000000000000000000000;
    wire [41:0] _38;
    wire [83:0] _40;
    wire [57:0] _41;
    wire [25:0] _36 = 26'b00000000000000000000000000;
    wire [83:0] _42;
    wire [15:0] _43;
    wire [31:0] _45;
    wire [15:0] _46;
    wire [15:0] _34;
    wire [15:0] _29 = 16'b0000000001100100;
    wire [41:0] _24 = 42'b000000000000000000000010100011110101110001;
    wire [25:0] _22 = 26'b00000000000000000000000000;
    wire [41:0] _23;
    wire [83:0] _25;
    wire [57:0] _26;
    wire [25:0] _21 = 26'b00000000000000000000000000;
    wire [83:0] _27;
    wire [15:0] _28;
    wire [31:0] _30;
    wire [15:0] _31;
    wire [15:0] _32;
    wire [15:0] _19 = 16'b0000000001100100;
    wire [15:0] _20;
    wire [15:0] _33;
    wire [15:0] _35;
    wire [15:0] _47;
    wire [15:0] _49;
    wire [15:0] _61;
    wire _63;
    wire [15:0] _69;
    wire _2;
    wire [15:0] _106;
    wire [15:0] _107;
    wire [15:0] _3;
    reg [15:0] _66;
    wire vdd = 1'b1;
    wire [15:0] _16 = 16'b0000000000000000;
    wire [15:0] _15 = 16'b0000000000000000;
    wire _6;
    wire [15:0] _137 = 16'b0000000000110010;
    wire [15:0] _133 = 16'b0000000001100100;
    wire [41:0] _128 = 42'b000000000000000000000010100011110101110001;
    wire [25:0] _126 = 26'b00000000000000000000000000;
    wire [41:0] _127;
    wire [83:0] _129;
    wire [57:0] _130;
    wire [25:0] _125 = 26'b00000000000000000000000000;
    wire [83:0] _131;
    wire [15:0] _132;
    wire [31:0] _134;
    wire [15:0] _135;
    wire [15:0] _123;
    wire [15:0] _118 = 16'b0000000001100100;
    wire [41:0] _113 = 42'b000000000000000000000010100011110101110001;
    wire [25:0] _111 = 26'b00000000000000000000000000;
    wire [41:0] _112;
    wire [83:0] _114;
    wire [57:0] _115;
    wire [25:0] _110 = 26'b00000000000000000000000000;
    wire [83:0] _116;
    wire [15:0] _117;
    wire [31:0] _119;
    wire [15:0] _120;
    wire [15:0] _8;
    wire [15:0] _121;
    wire [15:0] _108 = 16'b0000000001100100;
    wire [15:0] _109;
    wire [15:0] _122;
    wire _10;
    wire [15:0] _124;
    wire [15:0] _136;
    wire _12;
    wire [15:0] _138;
    wire [15:0] _13;
    reg [15:0] _18;

    /* logic */
    assign _102 = _49 == _62;
    assign _100 = _18 == _62;
    assign _101 = ~ _100;
    assign _103 = _101 & _102;
    assign _104 = _103 ? _67 : _62;
    assign _96 = _49 < _18;
    assign _92 = _49 == _62;
    assign _93 = ~ _92;
    assign _90 = _18 == _62;
    assign _91 = ~ _90;
    assign _94 = _91 & _93;
    assign _95 = _94 & _10;
    assign _97 = _95 & _96;
    assign _98 = _97 ? _67 : _62;
    assign _86 = _18 < _49;
    assign _84 = ~ _10;
    assign _81 = _49 == _62;
    assign _82 = ~ _81;
    assign _79 = _18 == _62;
    assign _80 = ~ _79;
    assign _83 = _80 & _82;
    assign _85 = _83 & _84;
    assign _87 = _85 & _86;
    assign _88 = _87 ? _67 : _62;
    assign _72 = { _71, _8 };
    assign _74 = _72 * _73;
    assign _75 = _74[83:26];
    assign _76 = { _70, _75 };
    assign _77 = _76[15:0];
    assign _78 = _66 + _77;
    assign _89 = _78 + _88;
    assign _99 = _89 + _98;
    assign _105 = _99 + _104;
    assign _68 = _66 + _67;
    assign _52 = { _51, _49 };
    assign _54 = _52 * _53;
    assign _55 = _54[83:26];
    assign _56 = { _50, _55 };
    assign _57 = _56[15:0];
    assign _59 = _57 * _58;
    assign _60 = _59[15:0];
    assign _38 = { _37, _35 };
    assign _40 = _38 * _39;
    assign _41 = _40[83:26];
    assign _42 = { _36, _41 };
    assign _43 = _42[15:0];
    assign _45 = _43 * _44;
    assign _46 = _45[15:0];
    assign _34 = _18 + _32;
    assign _23 = { _22, _8 };
    assign _25 = _23 * _24;
    assign _26 = _25[83:26];
    assign _27 = { _21, _26 };
    assign _28 = _27[15:0];
    assign _30 = _28 * _29;
    assign _31 = _30[15:0];
    assign _32 = _8 - _31;
    assign _20 = _18 + _19;
    assign _33 = _20 - _32;
    assign _35 = _10 ? _34 : _33;
    assign _47 = _35 - _46;
    assign _49 = _12 ? _48 : _47;
    assign _61 = _49 - _60;
    assign _63 = _61 == _62;
    assign _69 = _63 ? _68 : _66;
    assign _2 = part;
    assign _106 = _2 ? _105 : _69;
    assign _107 = _12 ? _62 : _106;
    assign _3 = _107;
    always @(posedge _6) begin
        _66 <= _3;
    end
    assign _6 = clock;
    assign _127 = { _126, _124 };
    assign _129 = _127 * _128;
    assign _130 = _129[83:26];
    assign _131 = { _125, _130 };
    assign _132 = _131[15:0];
    assign _134 = _132 * _133;
    assign _135 = _134[15:0];
    assign _123 = _18 + _121;
    assign _112 = { _111, _8 };
    assign _114 = _112 * _113;
    assign _115 = _114[83:26];
    assign _116 = { _110, _115 };
    assign _117 = _116[15:0];
    assign _119 = _117 * _118;
    assign _120 = _119[15:0];
    assign _8 = value;
    assign _121 = _8 - _120;
    assign _109 = _18 + _108;
    assign _122 = _109 - _121;
    assign _10 = positive;
    assign _124 = _10 ? _123 : _122;
    assign _136 = _124 - _135;
    assign _12 = reset;
    assign _138 = _12 ? _137 : _136;
    assign _13 = _138;
    always @(posedge _6) begin
        _18 <= _13;
    end

    /* aliases */

    /* output assignments */
    assign counter = _18;
    assign result = _66;

endmodule
